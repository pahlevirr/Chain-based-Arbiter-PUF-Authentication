clock_divider_inst : clock_divider PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig,
		locked	 => locked_sig
	);
